* D:\eSim_tut\files\clkdivider\clkdivider.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/22/23 10:12:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  rst GND pulse		
v2  clk GND pulse		
U5  rst clk Net-_U4-Pad1_ Net-_U4-Pad2_ adc_bridge_2		
U1  rst plot_v1		
U2  clk plot_v1		
U6  Net-_U4-Pad3_ clko dac_bridge_1		
U3  clko plot_v1		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ clkdivider		

.end
